covergroup foo;
    coverpoint x;
    some_name: coverpoint y;
endgroup
