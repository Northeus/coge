covergroup test1;
    coverpoint foo;
    coverpoint bar
    {
        bins a[] = 0;
        bins b[] = {1, 2, 3};
        bins c[] = {4, 5, 6};
    }
endgroup
